module main

fn main() {
	println(rgb(0, 0, 0).cmyk())
}
