module main

fn main() {
	println(hex(0x6789))
}
