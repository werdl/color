module color

pub fn d65() (f64, f64, f64) { // illuminus D65
	return 95.0455927, 100.0, 108.905775
}
