module main

fn main() {
	println(rgb(160,157,43).cielab())
}

